* First line is ignored

.global gnd vdd

*** SUBCIRCUIT NOR FROM CELL NOR{sch}
.SUBCKT NOR A AorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 AorB B gnd gnd NMOS L=0.4U W=2U
Mnmos@2 gnd A AorB gnd NMOS L=0.4U W=2U
Mpmos@1 net@112 B AorB vdd PMOS L=0.4U W=2U
Mpmos@2 vdd A net@112 vdd PMOS L=0.4U W=2U
.ENDS NOR
