*** SPICE deck for cell NOR{sch} from library nor2
*** Created on Fri Feb 16, 2024 23:07:43
*** Last revised on Mon Mar 04, 2024 22:07:12
*** Written on Mon Mar 04, 2024 22:17:48 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

.global gnd vdd

*** TOP LEVEL CELL: NOR{sch}
Mnmos@1 AorB B gnd gnd NMOS L=0.4U W=2U
Mnmos@2 gnd A AorB gnd NMOS L=0.4U W=2U
Mpmos@1 net@112 B AorB vdd PMOS L=0.4U W=2U
Mpmos@2 vdd A net@112 vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'NOR{sch}'
.measure tran tf trig v(AorB) val=4.5 fall=1 td=4ns targ v(AorB) val=0.5 fall=1
vb B 0 DC pwl 10n 0 20n 5 100n 5 110n 0
vdd vdd 0 DC 5 
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 140n 0 170n 0 180n 5
.measure tran tr trig v(AorB) val=0.5 rise=1 td=4ns targ v(AorB) val=4.5 rise=1
.tran 200n
.include C:\electric\C5_models.txt
.END
